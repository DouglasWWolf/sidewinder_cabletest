
//================================================================================================
//    Date         Version     Who  Changes
// -----------------------------------------------------------------------------------------------
// 03-Dec-2023     1.0.0       DWW  Initial creation
//================================================================================================
localparam VERSION_MAJOR = 1;
localparam VERSION_MINOR = 0;
localparam VERSION_BUILD = 0;
localparam VERSION_RCAND = 0;

localparam VERSION_DAY   = 9;
localparam VERSION_MONTH = 12;
localparam VERSION_YEAR  = 2023;
